library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity top_module_tb is
end top_module_tb

architecture Behavioral of top_module tb is
    component fila

